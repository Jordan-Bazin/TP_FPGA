library ieee ;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity chenillard is
	port (
		clk : in std_logic;
		rst : in std_logic;
		chen : out std_logic_vector(9 downto 0);
	);
end chenillard;

architecture behavioral of chenillard is

begin

end behavioral;
